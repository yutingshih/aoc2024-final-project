module controller (
    input rst,
    input clk,
    input enable,
    output finish,

    output [3:0] row_id, // X-Bus
    output [4:0] col_id, // Y-Bus PE id
);
    
endmodule