module top #(
    parameter  = ;
)(
    ports
);


    
endmodule